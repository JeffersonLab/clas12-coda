-- 
-- Si5345 Rev D Configuration Register Export Header File
-- 
-- This file represents a series of Skyworks Si5345 Rev D
-- register writes that can be performed to load a single configuration
-- on a device. It was created by a Skyworks ClockBuilder Pro
-- export tool.
-- 
-- Part:		                                       Si5345 Rev D
-- Design ID:                                          sPHX_GTM
-- Includes Pre/Post Download Control Register Writes: Yes
-- Created By:                                         ClockBuilder Pro v4.1 [2021-09-22]
-- Timestamp:                                          2021-10-25 14:42:06 GMT-04:00
-- 
-- A complete design report corresponding to this export is included at the end
-- of this header file.
-- 
-- 
-- signed int address; /* 16-bit register address */
-- signed char value; /* 8-bit register data */

-- Autogenerated on 2022-05-09 13:15:02.953620
-- by regmap_h2vhd.py

library ieee;
use ieee.std_logic_1164.all;

package si5345_register_pkg is
  type ROM_REC_T is record
      reg  : std_logic_vector(15 downto 0);
      data : std_logic_vector(7 downto 0);
  end record;
  type ROM_ARRAY_T is array (0 to 525) of ROM_REC_T;

  constant SI5345_ROM : ROM_ARRAY_T := ( 
-- Start configuration preamble */
    000 => (reg => x"0b24", data => x"c0"),
    001 => (reg => x"0b25", data => x"00"),
    002 => (reg => x"0540", data => x"01"),
-- End configuration preamble */
-- Delay 300 msec */
-- Delay is worst case time for device to complete any calibration */
-- that is running due to device state change previous to this script */
-- being processed. */
-- Start configuration registers */
    003 => (reg => x"0006", data => x"00"),
    004 => (reg => x"0007", data => x"00"),
    005 => (reg => x"0008", data => x"00"),
    006 => (reg => x"000b", data => x"68"),
    007 => (reg => x"0016", data => x"02"),
    008 => (reg => x"0017", data => x"dc"),
    009 => (reg => x"0018", data => x"ee"),
    010 => (reg => x"0019", data => x"dd"),
    011 => (reg => x"001a", data => x"df"),
    012 => (reg => x"002b", data => x"02"),
    013 => (reg => x"002c", data => x"01"),
    014 => (reg => x"002d", data => x"01"),
    015 => (reg => x"002e", data => x"35"),
    016 => (reg => x"002f", data => x"00"),
    017 => (reg => x"0030", data => x"00"),
    018 => (reg => x"0031", data => x"00"),
    019 => (reg => x"0032", data => x"00"),
    020 => (reg => x"0033", data => x"00"),
    021 => (reg => x"0034", data => x"00"),
    022 => (reg => x"0035", data => x"00"),
    023 => (reg => x"0036", data => x"35"),
    024 => (reg => x"0037", data => x"00"),
    025 => (reg => x"0038", data => x"00"),
    026 => (reg => x"0039", data => x"00"),
    027 => (reg => x"003a", data => x"00"),
    028 => (reg => x"003b", data => x"00"),
    029 => (reg => x"003c", data => x"00"),
    030 => (reg => x"003d", data => x"00"),
    031 => (reg => x"003f", data => x"11"),
    032 => (reg => x"0040", data => x"04"),
    033 => (reg => x"0041", data => x"0c"),
    034 => (reg => x"0042", data => x"00"),
    035 => (reg => x"0043", data => x"00"),
    036 => (reg => x"0044", data => x"00"),
    037 => (reg => x"0045", data => x"0c"),
    038 => (reg => x"0046", data => x"32"),
    039 => (reg => x"0047", data => x"00"),
    040 => (reg => x"0048", data => x"00"),
    041 => (reg => x"0049", data => x"00"),
    042 => (reg => x"004a", data => x"32"),
    043 => (reg => x"004b", data => x"00"),
    044 => (reg => x"004c", data => x"00"),
    045 => (reg => x"004d", data => x"00"),
    046 => (reg => x"004e", data => x"05"),
    047 => (reg => x"004f", data => x"00"),
    048 => (reg => x"0050", data => x"0f"),
    049 => (reg => x"0051", data => x"03"),
    050 => (reg => x"0052", data => x"00"),
    051 => (reg => x"0053", data => x"00"),
    052 => (reg => x"0054", data => x"00"),
    053 => (reg => x"0055", data => x"03"),
    054 => (reg => x"0056", data => x"00"),
    055 => (reg => x"0057", data => x"00"),
    056 => (reg => x"0058", data => x"00"),
    057 => (reg => x"0059", data => x"01"),
    058 => (reg => x"005a", data => x"55"),
    059 => (reg => x"005b", data => x"55"),
    060 => (reg => x"005c", data => x"d5"),
    061 => (reg => x"005d", data => x"00"),
    062 => (reg => x"005e", data => x"00"),
    063 => (reg => x"005f", data => x"00"),
    064 => (reg => x"0060", data => x"00"),
    065 => (reg => x"0061", data => x"00"),
    066 => (reg => x"0062", data => x"00"),
    067 => (reg => x"0063", data => x"00"),
    068 => (reg => x"0064", data => x"00"),
    069 => (reg => x"0065", data => x"00"),
    070 => (reg => x"0066", data => x"00"),
    071 => (reg => x"0067", data => x"00"),
    072 => (reg => x"0068", data => x"00"),
    073 => (reg => x"0069", data => x"00"),
    074 => (reg => x"0092", data => x"02"),
    075 => (reg => x"0093", data => x"a0"),
    076 => (reg => x"0095", data => x"00"),
    077 => (reg => x"0096", data => x"80"),
    078 => (reg => x"0098", data => x"60"),
    079 => (reg => x"009a", data => x"02"),
    080 => (reg => x"009b", data => x"60"),
    081 => (reg => x"009d", data => x"08"),
    082 => (reg => x"009e", data => x"40"),
    083 => (reg => x"00a0", data => x"20"),
    084 => (reg => x"00a2", data => x"00"),
    085 => (reg => x"00a9", data => x"6e"),
    086 => (reg => x"00aa", data => x"61"),
    087 => (reg => x"00ab", data => x"00"),
    088 => (reg => x"00ac", data => x"00"),
    089 => (reg => x"00e5", data => x"00"),
    090 => (reg => x"00ea", data => x"0a"),
    091 => (reg => x"00eb", data => x"60"),
    092 => (reg => x"00ec", data => x"00"),
    093 => (reg => x"00ed", data => x"00"),
    094 => (reg => x"0102", data => x"01"),
    095 => (reg => x"0108", data => x"01"),
    096 => (reg => x"0109", data => x"09"),
    097 => (reg => x"010a", data => x"3b"),
    098 => (reg => x"010b", data => x"28"),
    099 => (reg => x"010d", data => x"01"),
    100 => (reg => x"010e", data => x"09"),
    101 => (reg => x"010f", data => x"3b"),
    102 => (reg => x"0110", data => x"28"),
    103 => (reg => x"0112", data => x"01"),
    104 => (reg => x"0113", data => x"09"),
    105 => (reg => x"0114", data => x"3b"),
    106 => (reg => x"0115", data => x"28"),
    107 => (reg => x"0117", data => x"01"),
    108 => (reg => x"0118", data => x"09"),
    109 => (reg => x"0119", data => x"3b"),
    110 => (reg => x"011a", data => x"28"),
    111 => (reg => x"011c", data => x"01"),
    112 => (reg => x"011d", data => x"09"),
    113 => (reg => x"011e", data => x"3b"),
    114 => (reg => x"011f", data => x"28"),
    115 => (reg => x"0121", data => x"06"),
    116 => (reg => x"0122", data => x"09"),
    117 => (reg => x"0123", data => x"3b"),
    118 => (reg => x"0124", data => x"28"),
    119 => (reg => x"0126", data => x"01"),
    120 => (reg => x"0127", data => x"09"),
    121 => (reg => x"0128", data => x"3b"),
    122 => (reg => x"0129", data => x"28"),
    123 => (reg => x"012b", data => x"01"),
    124 => (reg => x"012c", data => x"09"),
    125 => (reg => x"012d", data => x"3b"),
    126 => (reg => x"012e", data => x"28"),
    127 => (reg => x"0130", data => x"01"),
    128 => (reg => x"0131", data => x"09"),
    129 => (reg => x"0132", data => x"3b"),
    130 => (reg => x"0133", data => x"28"),
    131 => (reg => x"013a", data => x"01"),
    132 => (reg => x"013b", data => x"09"),
    133 => (reg => x"013c", data => x"3b"),
    134 => (reg => x"013d", data => x"28"),
    135 => (reg => x"013f", data => x"00"),
    136 => (reg => x"0140", data => x"00"),
    137 => (reg => x"0141", data => x"40"),
    138 => (reg => x"0142", data => x"ff"),
    139 => (reg => x"0206", data => x"00"),
    140 => (reg => x"0208", data => x"14"),
    141 => (reg => x"0209", data => x"00"),
    142 => (reg => x"020a", data => x"00"),
    143 => (reg => x"020b", data => x"00"),
    144 => (reg => x"020c", data => x"00"),
    145 => (reg => x"020d", data => x"00"),
    146 => (reg => x"020e", data => x"01"),
    147 => (reg => x"020f", data => x"00"),
    148 => (reg => x"0210", data => x"00"),
    149 => (reg => x"0211", data => x"00"),
    150 => (reg => x"0212", data => x"00"),
    151 => (reg => x"0213", data => x"00"),
    152 => (reg => x"0214", data => x"00"),
    153 => (reg => x"0215", data => x"00"),
    154 => (reg => x"0216", data => x"00"),
    155 => (reg => x"0217", data => x"00"),
    156 => (reg => x"0218", data => x"00"),
    157 => (reg => x"0219", data => x"00"),
    158 => (reg => x"021a", data => x"00"),
    159 => (reg => x"021b", data => x"00"),
    160 => (reg => x"021c", data => x"00"),
    161 => (reg => x"021d", data => x"00"),
    162 => (reg => x"021e", data => x"00"),
    163 => (reg => x"021f", data => x"00"),
    164 => (reg => x"0220", data => x"00"),
    165 => (reg => x"0221", data => x"00"),
    166 => (reg => x"0222", data => x"00"),
    167 => (reg => x"0223", data => x"00"),
    168 => (reg => x"0224", data => x"00"),
    169 => (reg => x"0225", data => x"00"),
    170 => (reg => x"0226", data => x"00"),
    171 => (reg => x"0227", data => x"00"),
    172 => (reg => x"0228", data => x"00"),
    173 => (reg => x"0229", data => x"00"),
    174 => (reg => x"022a", data => x"00"),
    175 => (reg => x"022b", data => x"00"),
    176 => (reg => x"022c", data => x"00"),
    177 => (reg => x"022d", data => x"00"),
    178 => (reg => x"022e", data => x"00"),
    179 => (reg => x"022f", data => x"00"),
    180 => (reg => x"0231", data => x"0b"),
    181 => (reg => x"0232", data => x"0b"),
    182 => (reg => x"0233", data => x"0b"),
    183 => (reg => x"0234", data => x"0b"),
    184 => (reg => x"0235", data => x"00"),
    185 => (reg => x"0236", data => x"00"),
    186 => (reg => x"0237", data => x"00"),
    187 => (reg => x"0238", data => x"80"),
    188 => (reg => x"0239", data => x"89"),
    189 => (reg => x"023a", data => x"00"),
    190 => (reg => x"023b", data => x"00"),
    191 => (reg => x"023c", data => x"00"),
    192 => (reg => x"023d", data => x"00"),
    193 => (reg => x"023e", data => x"80"),
    194 => (reg => x"024a", data => x"00"),
    195 => (reg => x"024b", data => x"00"),
    196 => (reg => x"024c", data => x"00"),
    197 => (reg => x"024d", data => x"00"),
    198 => (reg => x"024e", data => x"00"),
    199 => (reg => x"024f", data => x"00"),
    200 => (reg => x"0250", data => x"00"),
    201 => (reg => x"0251", data => x"00"),
    202 => (reg => x"0252", data => x"00"),
    203 => (reg => x"0253", data => x"00"),
    204 => (reg => x"0254", data => x"00"),
    205 => (reg => x"0255", data => x"00"),
    206 => (reg => x"0256", data => x"00"),
    207 => (reg => x"0257", data => x"00"),
    208 => (reg => x"0258", data => x"00"),
    209 => (reg => x"0259", data => x"00"),
    210 => (reg => x"025a", data => x"00"),
    211 => (reg => x"025b", data => x"00"),
    212 => (reg => x"025c", data => x"00"),
    213 => (reg => x"025d", data => x"00"),
    214 => (reg => x"025e", data => x"00"),
    215 => (reg => x"025f", data => x"00"),
    216 => (reg => x"0260", data => x"00"),
    217 => (reg => x"0261", data => x"00"),
    218 => (reg => x"0262", data => x"00"),
    219 => (reg => x"0263", data => x"00"),
    220 => (reg => x"0264", data => x"00"),
    221 => (reg => x"0268", data => x"00"),
    222 => (reg => x"0269", data => x"00"),
    223 => (reg => x"026a", data => x"00"),
    224 => (reg => x"026b", data => x"73"),
    225 => (reg => x"026c", data => x"50"),
    226 => (reg => x"026d", data => x"48"),
    227 => (reg => x"026e", data => x"58"),
    228 => (reg => x"026f", data => x"5f"),
    229 => (reg => x"0270", data => x"47"),
    230 => (reg => x"0271", data => x"54"),
    231 => (reg => x"0272", data => x"4d"),
    232 => (reg => x"028a", data => x"00"),
    233 => (reg => x"028b", data => x"00"),
    234 => (reg => x"028c", data => x"00"),
    235 => (reg => x"028d", data => x"00"),
    236 => (reg => x"028e", data => x"00"),
    237 => (reg => x"028f", data => x"00"),
    238 => (reg => x"0290", data => x"00"),
    239 => (reg => x"0291", data => x"00"),
    240 => (reg => x"0294", data => x"b0"),
    241 => (reg => x"0296", data => x"02"),
    242 => (reg => x"0297", data => x"02"),
    243 => (reg => x"0299", data => x"02"),
    244 => (reg => x"029d", data => x"fa"),
    245 => (reg => x"029e", data => x"01"),
    246 => (reg => x"029f", data => x"00"),
    247 => (reg => x"02a9", data => x"cc"),
    248 => (reg => x"02aa", data => x"04"),
    249 => (reg => x"02ab", data => x"00"),
    250 => (reg => x"02b7", data => x"ff"),
    251 => (reg => x"0302", data => x"00"),
    252 => (reg => x"0303", data => x"00"),
    253 => (reg => x"0304", data => x"00"),
    254 => (reg => x"0305", data => x"80"),
    255 => (reg => x"0306", data => x"1b"),
    256 => (reg => x"0307", data => x"00"),
    257 => (reg => x"0308", data => x"00"),
    258 => (reg => x"0309", data => x"00"),
    259 => (reg => x"030a", data => x"00"),
    260 => (reg => x"030b", data => x"80"),
    261 => (reg => x"030c", data => x"00"),
    262 => (reg => x"030d", data => x"00"),
    263 => (reg => x"030e", data => x"00"),
    264 => (reg => x"030f", data => x"00"),
    265 => (reg => x"0310", data => x"00"),
    266 => (reg => x"0311", data => x"00"),
    267 => (reg => x"0312", data => x"00"),
    268 => (reg => x"0313", data => x"00"),
    269 => (reg => x"0314", data => x"00"),
    270 => (reg => x"0315", data => x"00"),
    271 => (reg => x"0316", data => x"00"),
    272 => (reg => x"0317", data => x"00"),
    273 => (reg => x"0318", data => x"00"),
    274 => (reg => x"0319", data => x"00"),
    275 => (reg => x"031a", data => x"00"),
    276 => (reg => x"031b", data => x"00"),
    277 => (reg => x"031c", data => x"00"),
    278 => (reg => x"031d", data => x"00"),
    279 => (reg => x"031e", data => x"00"),
    280 => (reg => x"031f", data => x"00"),
    281 => (reg => x"0320", data => x"00"),
    282 => (reg => x"0321", data => x"00"),
    283 => (reg => x"0322", data => x"00"),
    284 => (reg => x"0323", data => x"00"),
    285 => (reg => x"0324", data => x"00"),
    286 => (reg => x"0325", data => x"00"),
    287 => (reg => x"0326", data => x"00"),
    288 => (reg => x"0327", data => x"00"),
    289 => (reg => x"0328", data => x"00"),
    290 => (reg => x"0329", data => x"00"),
    291 => (reg => x"032a", data => x"00"),
    292 => (reg => x"032b", data => x"00"),
    293 => (reg => x"032c", data => x"00"),
    294 => (reg => x"032d", data => x"00"),
    295 => (reg => x"032e", data => x"00"),
    296 => (reg => x"032f", data => x"00"),
    297 => (reg => x"0330", data => x"00"),
    298 => (reg => x"0331", data => x"00"),
    299 => (reg => x"0332", data => x"00"),
    300 => (reg => x"0333", data => x"00"),
    301 => (reg => x"0334", data => x"00"),
    302 => (reg => x"0335", data => x"00"),
    303 => (reg => x"0336", data => x"00"),
    304 => (reg => x"0337", data => x"00"),
    305 => (reg => x"0338", data => x"00"),
    306 => (reg => x"0339", data => x"1f"),
    307 => (reg => x"033b", data => x"00"),
    308 => (reg => x"033c", data => x"00"),
    309 => (reg => x"033d", data => x"00"),
    310 => (reg => x"033e", data => x"00"),
    311 => (reg => x"033f", data => x"00"),
    312 => (reg => x"0340", data => x"00"),
    313 => (reg => x"0341", data => x"00"),
    314 => (reg => x"0342", data => x"00"),
    315 => (reg => x"0343", data => x"00"),
    316 => (reg => x"0344", data => x"00"),
    317 => (reg => x"0345", data => x"00"),
    318 => (reg => x"0346", data => x"00"),
    319 => (reg => x"0347", data => x"00"),
    320 => (reg => x"0348", data => x"00"),
    321 => (reg => x"0349", data => x"00"),
    322 => (reg => x"034a", data => x"00"),
    323 => (reg => x"034b", data => x"00"),
    324 => (reg => x"034c", data => x"00"),
    325 => (reg => x"034d", data => x"00"),
    326 => (reg => x"034e", data => x"00"),
    327 => (reg => x"034f", data => x"00"),
    328 => (reg => x"0350", data => x"00"),
    329 => (reg => x"0351", data => x"00"),
    330 => (reg => x"0352", data => x"00"),
    331 => (reg => x"0353", data => x"00"),
    332 => (reg => x"0354", data => x"00"),
    333 => (reg => x"0355", data => x"00"),
    334 => (reg => x"0356", data => x"00"),
    335 => (reg => x"0357", data => x"00"),
    336 => (reg => x"0358", data => x"00"),
    337 => (reg => x"0359", data => x"00"),
    338 => (reg => x"035a", data => x"00"),
    339 => (reg => x"035b", data => x"00"),
    340 => (reg => x"035c", data => x"00"),
    341 => (reg => x"035d", data => x"00"),
    342 => (reg => x"035e", data => x"00"),
    343 => (reg => x"035f", data => x"00"),
    344 => (reg => x"0360", data => x"00"),
    345 => (reg => x"0361", data => x"00"),
    346 => (reg => x"0362", data => x"00"),
    347 => (reg => x"0487", data => x"00"),
    348 => (reg => x"0508", data => x"13"),
    349 => (reg => x"0509", data => x"22"),
    350 => (reg => x"050a", data => x"0c"),
    351 => (reg => x"050b", data => x"0b"),
    352 => (reg => x"050c", data => x"07"),
    353 => (reg => x"050d", data => x"3f"),
    354 => (reg => x"050e", data => x"16"),
    355 => (reg => x"050f", data => x"2a"),
    356 => (reg => x"0510", data => x"09"),
    357 => (reg => x"0511", data => x"08"),
    358 => (reg => x"0512", data => x"07"),
    359 => (reg => x"0513", data => x"3f"),
    360 => (reg => x"0515", data => x"00"),
    361 => (reg => x"0516", data => x"00"),
    362 => (reg => x"0517", data => x"00"),
    363 => (reg => x"0518", data => x"00"),
    364 => (reg => x"0519", data => x"94"),
    365 => (reg => x"051a", data => x"02"),
    366 => (reg => x"051b", data => x"00"),
    367 => (reg => x"051c", data => x"00"),
    368 => (reg => x"051d", data => x"00"),
    369 => (reg => x"051e", data => x"00"),
    370 => (reg => x"051f", data => x"80"),
    371 => (reg => x"0521", data => x"2b"),
    372 => (reg => x"052a", data => x"01"),
    373 => (reg => x"052b", data => x"01"),
    374 => (reg => x"052c", data => x"87"),
    375 => (reg => x"052d", data => x"03"),
    376 => (reg => x"052e", data => x"19"),
    377 => (reg => x"052f", data => x"19"),
    378 => (reg => x"0531", data => x"00"),
    379 => (reg => x"0532", data => x"42"),
    380 => (reg => x"0533", data => x"03"),
    381 => (reg => x"0534", data => x"00"),
    382 => (reg => x"0535", data => x"00"),
    383 => (reg => x"0536", data => x"00"),
    384 => (reg => x"0537", data => x"00"),
    385 => (reg => x"0538", data => x"00"),
    386 => (reg => x"0539", data => x"00"),
    387 => (reg => x"053a", data => x"02"),
    388 => (reg => x"053b", data => x"03"),
    389 => (reg => x"053c", data => x"00"),
    390 => (reg => x"053d", data => x"11"),
    391 => (reg => x"053e", data => x"06"),
    392 => (reg => x"0589", data => x"0d"),
    393 => (reg => x"058a", data => x"00"),
    394 => (reg => x"059b", data => x"f8"),
    395 => (reg => x"059d", data => x"13"),
    396 => (reg => x"059e", data => x"24"),
    397 => (reg => x"059f", data => x"0c"),
    398 => (reg => x"05a0", data => x"0b"),
    399 => (reg => x"05a1", data => x"07"),
    400 => (reg => x"05a2", data => x"3f"),
    401 => (reg => x"05a6", data => x"03"),
    402 => (reg => x"0802", data => x"35"),
    403 => (reg => x"0803", data => x"05"),
    404 => (reg => x"0804", data => x"00"),
    405 => (reg => x"0805", data => x"00"),
    406 => (reg => x"0806", data => x"00"),
    407 => (reg => x"0807", data => x"00"),
    408 => (reg => x"0808", data => x"00"),
    409 => (reg => x"0809", data => x"00"),
    410 => (reg => x"080a", data => x"00"),
    411 => (reg => x"080b", data => x"00"),
    412 => (reg => x"080c", data => x"00"),
    413 => (reg => x"080d", data => x"00"),
    414 => (reg => x"080e", data => x"00"),
    415 => (reg => x"080f", data => x"00"),
    416 => (reg => x"0810", data => x"00"),
    417 => (reg => x"0811", data => x"00"),
    418 => (reg => x"0812", data => x"00"),
    419 => (reg => x"0813", data => x"00"),
    420 => (reg => x"0814", data => x"00"),
    421 => (reg => x"0815", data => x"00"),
    422 => (reg => x"0816", data => x"00"),
    423 => (reg => x"0817", data => x"00"),
    424 => (reg => x"0818", data => x"00"),
    425 => (reg => x"0819", data => x"00"),
    426 => (reg => x"081a", data => x"00"),
    427 => (reg => x"081b", data => x"00"),
    428 => (reg => x"081c", data => x"00"),
    429 => (reg => x"081d", data => x"00"),
    430 => (reg => x"081e", data => x"00"),
    431 => (reg => x"081f", data => x"00"),
    432 => (reg => x"0820", data => x"00"),
    433 => (reg => x"0821", data => x"00"),
    434 => (reg => x"0822", data => x"00"),
    435 => (reg => x"0823", data => x"00"),
    436 => (reg => x"0824", data => x"00"),
    437 => (reg => x"0825", data => x"00"),
    438 => (reg => x"0826", data => x"00"),
    439 => (reg => x"0827", data => x"00"),
    440 => (reg => x"0828", data => x"00"),
    441 => (reg => x"0829", data => x"00"),
    442 => (reg => x"082a", data => x"00"),
    443 => (reg => x"082b", data => x"00"),
    444 => (reg => x"082c", data => x"00"),
    445 => (reg => x"082d", data => x"00"),
    446 => (reg => x"082e", data => x"00"),
    447 => (reg => x"082f", data => x"00"),
    448 => (reg => x"0830", data => x"00"),
    449 => (reg => x"0831", data => x"00"),
    450 => (reg => x"0832", data => x"00"),
    451 => (reg => x"0833", data => x"00"),
    452 => (reg => x"0834", data => x"00"),
    453 => (reg => x"0835", data => x"00"),
    454 => (reg => x"0836", data => x"00"),
    455 => (reg => x"0837", data => x"00"),
    456 => (reg => x"0838", data => x"00"),
    457 => (reg => x"0839", data => x"00"),
    458 => (reg => x"083a", data => x"00"),
    459 => (reg => x"083b", data => x"00"),
    460 => (reg => x"083c", data => x"00"),
    461 => (reg => x"083d", data => x"00"),
    462 => (reg => x"083e", data => x"00"),
    463 => (reg => x"083f", data => x"00"),
    464 => (reg => x"0840", data => x"00"),
    465 => (reg => x"0841", data => x"00"),
    466 => (reg => x"0842", data => x"00"),
    467 => (reg => x"0843", data => x"00"),
    468 => (reg => x"0844", data => x"00"),
    469 => (reg => x"0845", data => x"00"),
    470 => (reg => x"0846", data => x"00"),
    471 => (reg => x"0847", data => x"00"),
    472 => (reg => x"0848", data => x"00"),
    473 => (reg => x"0849", data => x"00"),
    474 => (reg => x"084a", data => x"00"),
    475 => (reg => x"084b", data => x"00"),
    476 => (reg => x"084c", data => x"00"),
    477 => (reg => x"084d", data => x"00"),
    478 => (reg => x"084e", data => x"00"),
    479 => (reg => x"084f", data => x"00"),
    480 => (reg => x"0850", data => x"00"),
    481 => (reg => x"0851", data => x"00"),
    482 => (reg => x"0852", data => x"00"),
    483 => (reg => x"0853", data => x"00"),
    484 => (reg => x"0854", data => x"00"),
    485 => (reg => x"0855", data => x"00"),
    486 => (reg => x"0856", data => x"00"),
    487 => (reg => x"0857", data => x"00"),
    488 => (reg => x"0858", data => x"00"),
    489 => (reg => x"0859", data => x"00"),
    490 => (reg => x"085a", data => x"00"),
    491 => (reg => x"085b", data => x"00"),
    492 => (reg => x"085c", data => x"00"),
    493 => (reg => x"085d", data => x"00"),
    494 => (reg => x"085e", data => x"00"),
    495 => (reg => x"085f", data => x"00"),
    496 => (reg => x"0860", data => x"00"),
    497 => (reg => x"0861", data => x"00"),
    498 => (reg => x"090e", data => x"02"),
    499 => (reg => x"0943", data => x"00"),
    500 => (reg => x"0949", data => x"01"),
    501 => (reg => x"094a", data => x"01"),
    502 => (reg => x"094e", data => x"49"),
    503 => (reg => x"094f", data => x"02"),
    504 => (reg => x"095e", data => x"00"),
    505 => (reg => x"0a02", data => x"00"),
    506 => (reg => x"0a03", data => x"01"),
    507 => (reg => x"0a04", data => x"01"),
    508 => (reg => x"0a05", data => x"01"),
    509 => (reg => x"0a14", data => x"00"),
    510 => (reg => x"0a1a", data => x"00"),
    511 => (reg => x"0a20", data => x"00"),
    512 => (reg => x"0a26", data => x"00"),
    513 => (reg => x"0a2c", data => x"00"),
    514 => (reg => x"0b44", data => x"2f"),
    515 => (reg => x"0b46", data => x"00"),
    516 => (reg => x"0b47", data => x"0e"),
    517 => (reg => x"0b48", data => x"0e"),
    518 => (reg => x"0b4a", data => x"1e"),
    519 => (reg => x"0b57", data => x"0e"),
    520 => (reg => x"0b58", data => x"01"),
-- End configuration registers */
-- Start configuration postamble */
    521 => (reg => x"0514", data => x"01"),
    522 => (reg => x"001c", data => x"01"),
    523 => (reg => x"0540", data => x"00"),
    524 => (reg => x"0b24", data => x"c3"),
-- End configuration postamble */
    525 => (reg => x"0b25", data => x"02")
  );
-- 
-- Design Report
-- 
-- Overview
-- ========
-- Part:               Si5345ABCD Rev D
-- Design ID:          sPHX_GTM
-- Created By:         ClockBuilder Pro v4.1 [2021-09-22]
-- Timestamp:          2021-10-25 14:42:06 GMT-04:00
-- 
-- Design Rule Check
-- =================
-- Errors:
-- - No errors
-- 
-- Warnings:
-- - No warnings
-- 
-- Device Grade
-- ============
-- Maximum Output Frequency: 120 MHz
-- Frequency Synthesis Mode: Integer
-- Frequency Plan Grade:     D
-- Minimum Base OPN:         Si5345D*
-- 
-- Base       Output Clock         Supported Frequency Synthesis Modes
-- OPN Grade  Frequency Range      (Typical Jitter)
-- ---------  -------------------  --------------------------------------------
-- Si5345A    100 Hz to 1.028 GHz  Integer (< 100 fs) and fractional (< 150 fs)
-- Si5345B    100 Hz to 350 MHz    "
-- Si5345C    100 Hz to 1.028 GHz  Integer only (< 100 fs)
-- Si5345D*   100 Hz to 350 MHz    "
-- 
-- * Based on your calculated frequency plan, a Si5345D grade device is
-- sufficient for your design. For more in-system configuration flexibility
-- (higher frequencies and/or to enable fractional synthesis), consider
-- selecting device grade Si5345A when specifying an ordering part number (OPN)
-- for your application. See the datasheet Ordering Guide for more information.
-- 
-- Design
-- ======
-- Host Interface:
-- I/O Power Supply: VDD (Core)
-- SPI Mode: 4-Wire
-- I2C Address Range: 104d to 107d / 0x68 to 0x6B (selected via A0/A1 pins)
-- 
-- XA/XB:
-- 48 MHz (XTAL - Crystal)
-- 
-- Inputs:
-- IN0: 40 MHz
-- Standard
-- IN1: Unused
-- IN2: Unused
-- IN3: Unused
-- 
-- Outputs:
-- OUT0: Unused
-- OUT1: Unused
-- OUT2: Unused
-- OUT3: Unused
-- OUT4: Unused
-- OUT5: 120 MHz
-- Enabled, LVDS 2.5 V
-- OUT6: Unused
-- OUT7: Unused
-- OUT8: Unused
-- OUT9: Unused
-- 
-- Frequency Plan
-- ==============
-- Priority: maximize the number of low jitter outputs
-- 
-- Fvco = 13.2 GHz
-- Fpfd = 2 MHz
-- Fms0 = 240 MHz
-- 
-- P dividers:
-- P0  = 20
-- P1  = Unused
-- P2  = Unused
-- P3  = Unused
-- Pxaxb = 1
-- 
-- MXAXB = 275
-- M = 1320
-- N dividers:
-- N0:
-- Value: 55
-- OUT5: 120 MHz
-- N1:
-- Unused
-- N2:
-- Unused
-- N3:
-- Unused
-- N4:
-- Unused
-- 
-- R dividers:
-- R0 = Unused
-- R1 = Unused
-- R2 = Unused
-- R3 = Unused
-- R4 = Unused
-- R5 = 2
-- R6 = Unused
-- R7 = Unused
-- R8 = Unused
-- R9 = Unused
-- 
-- Nominal Bandwidth:
-- Desired: 100.000 Hz
-- Actual:  92.196 Hz
-- Coefficients:
-- BW0:  19
-- BW1:  34
-- BW2:  12
-- BW3:  11
-- BW4:  7
-- BW5:  63
-- Fastlock Bandwidth:
-- Desired: 1.000 kHz
-- Actual:  738.336 Hz
-- Coefficients:
-- BW0:  22
-- BW1:  42
-- BW2:  9
-- BW3:  8
-- BW4:  7
-- BW5:  63
-- Holdover Bandwidth:
-- N/A (Ramped Exit from Holdover)
-- 
-- Dividers listed above show effective values. These values are translated to register settings by ClockBuilder Pro. For the actual register values, see below. Refer to the Family Reference Manual for information on registers related to frequency plan.
-- 
-- Digitally Controlled Oscillator (DCO)
-- =====================================
-- Mode: Register Direct Write
-- 
-- N0: DCO Disabled
-- 
-- N1: DCO Disabled
-- 
-- N2: DCO Disabled
-- 
-- N3: DCO Disabled
-- 
-- N4: DCO Disabled
-- 
-- Estimated Power & Junction Temperature
-- ======================================
-- Assumptions:
-- 
-- Revision: D
-- VDD:      1.8 V
-- Ta:       25 �C
-- Theta-JA: 18.3 �C/W
-- Airflow:  2 m/s
-- 
-- Total Power: 602 mW, On Chip Power: 596 mW, Tj: 36 �C
-- 
-- Frequency  Format   Voltage   Current     Power
-- ---------  ------  --------  --------  --------
-- VDD                           1.8 V  102.2 mA    184 mW
-- VDDA                          3.3 V  114.8 mA    379 mW
-- VDDO0      Unused
-- VDDO1      Unused
-- VDDO2      Unused
-- VDDO3      Unused
-- VDDO4      Unused
-- VDDO5     120 MHz  LVDS       2.5 V   15.6 mA     39 mW
-- VDDO6      Unused
-- VDDO7      Unused
-- VDDO8      Unused
-- VDDO9      Unused
-- --------  --------
-- Total  232.5 mA    602 mW
-- 
-- Note:
-- 
-- -Tj is junction temperature. Tj must be less than 125 �C (on Si5345 Revision D) for device to comply with datasheet specifications. Tj = Ta + Theta_JA*On_Chip_Power.
-- -Overall power includes on-chip power dissipation and adds differential load power dissipation to estimate total power requirements.
-- -Above are estimates only: power and temperature should be measured on your PCB.
-- -Selection of appropriate Theta-JA is required for most accurate estimate. Ideally, select 'User Specified Theta-JA' and enter a Theta-JA value based on the thermal properties of your PCB.
-- 
-- Settings
-- ========
-- 
-- Location      Setting Name                Decimal Value      Hex Value
-- ------------  --------------------------  -----------------  -----------------
-- 0x0006[23:0]  TOOL_VERSION                0                  0x000000
-- 0x000B[6:0]   I2C_ADDR                    104                0x68
-- 0x0016[1]     LOL_ON_HOLD                 1                  0x1
-- 0x0017[0]     SYSINCAL_INTR_MSK           0                  0x0
-- 0x0017[1]     LOSXAXB_INTR_MSK            0                  0x0
-- 0x0017[5]     SMB_TMOUT_INTR_MSK          0                  0x0
-- 0x0018[3:0]   LOS_INTR_MSK                14                 0xE
-- 0x0018[7:4]   OOF_INTR_MSK                14                 0xE
-- 0x0019[1]     LOL_INTR_MSK                0                  0x0
-- 0x0019[5]     HOLD_INTR_MSK               0                  0x0
-- 0x001A[5]     CAL_INTR_MSK                0                  0x0
-- 0x002B[3]     SPI_3WIRE                   0                  0x0
-- 0x002B[5]     AUTO_NDIV_UPDATE            0                  0x0
-- 0x002C[3:0]   LOS_EN                      1                  0x1
-- 0x002C[4]     LOSXAXB_DIS                 0                  0x0
-- 0x002D[1:0]   LOS0_VAL_TIME               1                  0x1
-- 0x002D[3:2]   LOS1_VAL_TIME               0                  0x0
-- 0x002D[5:4]   LOS2_VAL_TIME               0                  0x0
-- 0x002D[7:6]   LOS3_VAL_TIME               0                  0x0
-- 0x002E[15:0]  LOS0_TRG_THR                53                 0x0035
-- 0x0030[15:0]  LOS1_TRG_THR                0                  0x0000
-- 0x0032[15:0]  LOS2_TRG_THR                0                  0x0000
-- 0x0034[15:0]  LOS3_TRG_THR                0                  0x0000
-- 0x0036[15:0]  LOS0_CLR_THR                53                 0x0035
-- 0x0038[15:0]  LOS1_CLR_THR                0                  0x0000
-- 0x003A[15:0]  LOS2_CLR_THR                0                  0x0000
-- 0x003C[15:0]  LOS3_CLR_THR                0                  0x0000
-- 0x003F[3:0]   OOF_EN                      1                  0x1
-- 0x003F[7:4]   FAST_OOF_EN                 1                  0x1
-- 0x0040[2:0]   OOF_REF_SEL                 4                  0x4
-- 0x0041[4:0]   OOF0_DIV_SEL                12                 0x0C
-- 0x0042[4:0]   OOF1_DIV_SEL                0                  0x00
-- 0x0043[4:0]   OOF2_DIV_SEL                0                  0x00
-- 0x0044[4:0]   OOF3_DIV_SEL                0                  0x00
-- 0x0045[4:0]   OOFXO_DIV_SEL               12                 0x0C
-- 0x0046[7:0]   OOF0_SET_THR                50                 0x32
-- 0x0047[7:0]   OOF1_SET_THR                0                  0x00
-- 0x0048[7:0]   OOF2_SET_THR                0                  0x00
-- 0x0049[7:0]   OOF3_SET_THR                0                  0x00
-- 0x004A[7:0]   OOF0_CLR_THR                50                 0x32
-- 0x004B[7:0]   OOF1_CLR_THR                0                  0x00
-- 0x004C[7:0]   OOF2_CLR_THR                0                  0x00
-- 0x004D[7:0]   OOF3_CLR_THR                0                  0x00
-- 0x004E[2:0]   OOF0_DETWIN_SEL             5                  0x5
-- 0x004E[6:4]   OOF1_DETWIN_SEL             0                  0x0
-- 0x004F[2:0]   OOF2_DETWIN_SEL             0                  0x0
-- 0x004F[6:4]   OOF3_DETWIN_SEL             0                  0x0
-- 0x0050[3:0]   OOF_ON_LOS                  15                 0xF
-- 0x0051[3:0]   FAST_OOF0_SET_THR           3                  0x3
-- 0x0052[3:0]   FAST_OOF1_SET_THR           0                  0x0
-- 0x0053[3:0]   FAST_OOF2_SET_THR           0                  0x0
-- 0x0054[3:0]   FAST_OOF3_SET_THR           0                  0x0
-- 0x0055[3:0]   FAST_OOF0_CLR_THR           3                  0x3
-- 0x0056[3:0]   FAST_OOF1_CLR_THR           0                  0x0
-- 0x0057[3:0]   FAST_OOF2_CLR_THR           0                  0x0
-- 0x0058[3:0]   FAST_OOF3_CLR_THR           0                  0x0
-- 0x0059[1:0]   FAST_OOF0_DETWIN_SEL        1                  0x1
-- 0x0059[3:2]   FAST_OOF1_DETWIN_SEL        0                  0x0
-- 0x0059[5:4]   FAST_OOF2_DETWIN_SEL        0                  0x0
-- 0x0059[7:6]   FAST_OOF3_DETWIN_SEL        0                  0x0
-- 0x005A[25:0]  OOF0_RATIO_REF              13981013           0x0D55555
-- 0x005E[25:0]  OOF1_RATIO_REF              0                  0x0000000
-- 0x0062[25:0]  OOF2_RATIO_REF              0                  0x0000000
-- 0x0066[25:0]  OOF3_RATIO_REF              0                  0x0000000
-- 0x0092[1]     LOL_FST_EN                  1                  0x1
-- 0x0093[7:4]   LOL_FST_DETWIN_SEL          10                 0xA
-- 0x0095[3:2]   LOL_FST_VALWIN_SEL          0                  0x0
-- 0x0096[7:4]   LOL_FST_SET_THR_SEL         8                  0x8
-- 0x0098[7:4]   LOL_FST_CLR_THR_SEL         6                  0x6
-- 0x009A[1]     LOL_SLOW_EN_PLL             1                  0x1
-- 0x009B[7:4]   LOL_SLW_DETWIN_SEL          6                  0x6
-- 0x009D[3:2]   LOL_SLW_VALWIN_SEL          2                  0x2
-- 0x009E[7:4]   LOL_SLW_SET_THR             4                  0x4
-- 0x00A0[7:4]   LOL_SLW_CLR_THR             2                  0x2
-- 0x00A2[1]     LOL_TIMER_EN                0                  0x0
-- 0x00A9[28:0]  LOL_CLR_DELAY_DIV256        24942              0x0000616E
-- 0x00E5[0]     FASTLOCK_EXTEND_MASTER_DIS  0                  0x0
-- 0x00E5[5]     FASTLOCK_EXTEND_EN          0                  0x0
-- 0x00EA[28:0]  FASTLOCK_EXTEND             24586              0x0000600A
-- 0x0102[0]     OUTALL_DISABLE_LOW          1                  0x1
-- 0x0108[0]     OUT0_PDN                    1                  0x1
-- 0x0108[1]     OUT0_OE                     0                  0x0
-- 0x0108[2]     OUT0_RDIV_FORCE2            0                  0x0
-- 0x0109[2:0]   OUT0_FORMAT                 1                  0x1
-- 0x0109[3]     OUT0_SYNC_EN                1                  0x1
-- 0x0109[5:4]   OUT0_DIS_STATE              0                  0x0
-- 0x0109[7:6]   OUT0_CMOS_DRV               0                  0x0
-- 0x010A[3:0]   OUT0_CM                     11                 0xB
-- 0x010A[6:4]   OUT0_AMPL                   3                  0x3
-- 0x010B[2:0]   OUT0_MUX_SEL                0                  0x0
-- 0x010B[5:4]   OUT0_VDD_SEL                2                  0x2
-- 0x010B[3]     OUT0_VDD_SEL_EN             1                  0x1
-- 0x010B[7:6]   OUT0_INV                    0                  0x0
-- 0x010D[0]     OUT1_PDN                    1                  0x1
-- 0x010D[1]     OUT1_OE                     0                  0x0
-- 0x010D[2]     OUT1_RDIV_FORCE2            0                  0x0
-- 0x010E[2:0]   OUT1_FORMAT                 1                  0x1
-- 0x010E[3]     OUT1_SYNC_EN                1                  0x1
-- 0x010E[5:4]   OUT1_DIS_STATE              0                  0x0
-- 0x010E[7:6]   OUT1_CMOS_DRV               0                  0x0
-- 0x010F[3:0]   OUT1_CM                     11                 0xB
-- 0x010F[6:4]   OUT1_AMPL                   3                  0x3
-- 0x0110[2:0]   OUT1_MUX_SEL                0                  0x0
-- 0x0110[5:4]   OUT1_VDD_SEL                2                  0x2
-- 0x0110[3]     OUT1_VDD_SEL_EN             1                  0x1
-- 0x0110[7:6]   OUT1_INV                    0                  0x0
-- 0x0112[0]     OUT2_PDN                    1                  0x1
-- 0x0112[1]     OUT2_OE                     0                  0x0
-- 0x0112[2]     OUT2_RDIV_FORCE2            0                  0x0
-- 0x0113[2:0]   OUT2_FORMAT                 1                  0x1
-- 0x0113[3]     OUT2_SYNC_EN                1                  0x1
-- 0x0113[5:4]   OUT2_DIS_STATE              0                  0x0
-- 0x0113[7:6]   OUT2_CMOS_DRV               0                  0x0
-- 0x0114[3:0]   OUT2_CM                     11                 0xB
-- 0x0114[6:4]   OUT2_AMPL                   3                  0x3
-- 0x0115[2:0]   OUT2_MUX_SEL                0                  0x0
-- 0x0115[5:4]   OUT2_VDD_SEL                2                  0x2
-- 0x0115[3]     OUT2_VDD_SEL_EN             1                  0x1
-- 0x0115[7:6]   OUT2_INV                    0                  0x0
-- 0x0117[0]     OUT3_PDN                    1                  0x1
-- 0x0117[1]     OUT3_OE                     0                  0x0
-- 0x0117[2]     OUT3_RDIV_FORCE2            0                  0x0
-- 0x0118[2:0]   OUT3_FORMAT                 1                  0x1
-- 0x0118[3]     OUT3_SYNC_EN                1                  0x1
-- 0x0118[5:4]   OUT3_DIS_STATE              0                  0x0
-- 0x0118[7:6]   OUT3_CMOS_DRV               0                  0x0
-- 0x0119[3:0]   OUT3_CM                     11                 0xB
-- 0x0119[6:4]   OUT3_AMPL                   3                  0x3
-- 0x011A[2:0]   OUT3_MUX_SEL                0                  0x0
-- 0x011A[5:4]   OUT3_VDD_SEL                2                  0x2
-- 0x011A[3]     OUT3_VDD_SEL_EN             1                  0x1
-- 0x011A[7:6]   OUT3_INV                    0                  0x0
-- 0x011C[0]     OUT4_PDN                    1                  0x1
-- 0x011C[1]     OUT4_OE                     0                  0x0
-- 0x011C[2]     OUT4_RDIV_FORCE2            0                  0x0
-- 0x011D[2:0]   OUT4_FORMAT                 1                  0x1
-- 0x011D[3]     OUT4_SYNC_EN                1                  0x1
-- 0x011D[5:4]   OUT4_DIS_STATE              0                  0x0
-- 0x011D[7:6]   OUT4_CMOS_DRV               0                  0x0
-- 0x011E[3:0]   OUT4_CM                     11                 0xB
-- 0x011E[6:4]   OUT4_AMPL                   3                  0x3
-- 0x011F[2:0]   OUT4_MUX_SEL                0                  0x0
-- 0x011F[5:4]   OUT4_VDD_SEL                2                  0x2
-- 0x011F[3]     OUT4_VDD_SEL_EN             1                  0x1
-- 0x011F[7:6]   OUT4_INV                    0                  0x0
-- 0x0121[0]     OUT5_PDN                    0                  0x0
-- 0x0121[1]     OUT5_OE                     1                  0x1
-- 0x0121[2]     OUT5_RDIV_FORCE2            1                  0x1
-- 0x0122[2:0]   OUT5_FORMAT                 1                  0x1
-- 0x0122[3]     OUT5_SYNC_EN                1                  0x1
-- 0x0122[5:4]   OUT5_DIS_STATE              0                  0x0
-- 0x0122[7:6]   OUT5_CMOS_DRV               0                  0x0
-- 0x0123[3:0]   OUT5_CM                     11                 0xB
-- 0x0123[6:4]   OUT5_AMPL                   3                  0x3
-- 0x0124[2:0]   OUT5_MUX_SEL                0                  0x0
-- 0x0124[5:4]   OUT5_VDD_SEL                2                  0x2
-- 0x0124[3]     OUT5_VDD_SEL_EN             1                  0x1
-- 0x0124[7:6]   OUT5_INV                    0                  0x0
-- 0x0126[0]     OUT6_PDN                    1                  0x1
-- 0x0126[1]     OUT6_OE                     0                  0x0
-- 0x0126[2]     OUT6_RDIV_FORCE2            0                  0x0
-- 0x0127[2:0]   OUT6_FORMAT                 1                  0x1
-- 0x0127[3]     OUT6_SYNC_EN                1                  0x1
-- 0x0127[5:4]   OUT6_DIS_STATE              0                  0x0
-- 0x0127[7:6]   OUT6_CMOS_DRV               0                  0x0
-- 0x0128[3:0]   OUT6_CM                     11                 0xB
-- 0x0128[6:4]   OUT6_AMPL                   3                  0x3
-- 0x0129[2:0]   OUT6_MUX_SEL                0                  0x0
-- 0x0129[5:4]   OUT6_VDD_SEL                2                  0x2
-- 0x0129[3]     OUT6_VDD_SEL_EN             1                  0x1
-- 0x0129[7:6]   OUT6_INV                    0                  0x0
-- 0x012B[0]     OUT7_PDN                    1                  0x1
-- 0x012B[1]     OUT7_OE                     0                  0x0
-- 0x012B[2]     OUT7_RDIV_FORCE2            0                  0x0
-- 0x012C[2:0]   OUT7_FORMAT                 1                  0x1
-- 0x012C[3]     OUT7_SYNC_EN                1                  0x1
-- 0x012C[5:4]   OUT7_DIS_STATE              0                  0x0
-- 0x012C[7:6]   OUT7_CMOS_DRV               0                  0x0
-- 0x012D[3:0]   OUT7_CM                     11                 0xB
-- 0x012D[6:4]   OUT7_AMPL                   3                  0x3
-- 0x012E[2:0]   OUT7_MUX_SEL                0                  0x0
-- 0x012E[5:4]   OUT7_VDD_SEL                2                  0x2
-- 0x012E[3]     OUT7_VDD_SEL_EN             1                  0x1
-- 0x012E[7:6]   OUT7_INV                    0                  0x0
-- 0x0130[0]     OUT8_PDN                    1                  0x1
-- 0x0130[1]     OUT8_OE                     0                  0x0
-- 0x0130[2]     OUT8_RDIV_FORCE2            0                  0x0
-- 0x0131[2:0]   OUT8_FORMAT                 1                  0x1
-- 0x0131[3]     OUT8_SYNC_EN                1                  0x1
-- 0x0131[5:4]   OUT8_DIS_STATE              0                  0x0
-- 0x0131[7:6]   OUT8_CMOS_DRV               0                  0x0
-- 0x0132[3:0]   OUT8_CM                     11                 0xB
-- 0x0132[6:4]   OUT8_AMPL                   3                  0x3
-- 0x0133[2:0]   OUT8_MUX_SEL                0                  0x0
-- 0x0133[5:4]   OUT8_VDD_SEL                2                  0x2
-- 0x0133[3]     OUT8_VDD_SEL_EN             1                  0x1
-- 0x0133[7:6]   OUT8_INV                    0                  0x0
-- 0x013A[0]     OUT9_PDN                    1                  0x1
-- 0x013A[1]     OUT9_OE                     0                  0x0
-- 0x013A[2]     OUT9_RDIV_FORCE2            0                  0x0
-- 0x013B[2:0]   OUT9_FORMAT                 1                  0x1
-- 0x013B[3]     OUT9_SYNC_EN                1                  0x1
-- 0x013B[5:4]   OUT9_DIS_STATE              0                  0x0
-- 0x013B[7:6]   OUT9_CMOS_DRV               0                  0x0
-- 0x013C[3:0]   OUT9_CM                     11                 0xB
-- 0x013C[6:4]   OUT9_AMPL                   3                  0x3
-- 0x013D[2:0]   OUT9_MUX_SEL                0                  0x0
-- 0x013D[5:4]   OUT9_VDD_SEL                2                  0x2
-- 0x013D[3]     OUT9_VDD_SEL_EN             1                  0x1
-- 0x013D[7:6]   OUT9_INV                    0                  0x0
-- 0x013F[11:0]  OUTX_ALWAYS_ON              0                  0x000
-- 0x0141[1]     OUT_DIS_MSK                 0                  0x0
-- 0x0141[5]     OUT_DIS_LOL_MSK             0                  0x0
-- 0x0141[6]     OUT_DIS_LOSXAXB_MSK         1                  0x1
-- 0x0141[7]     OUT_DIS_MSK_LOS_PFD         0                  0x0
-- 0x0142[1]     OUT_DIS_MSK_LOL             1                  0x1
-- 0x0142[5]     OUT_DIS_MSK_HOLD            1                  0x1
-- 0x0206[1:0]   PXAXB                       0                  0x0
-- 0x0208[47:0]  P0_NUM                      20                 0x000000000014
-- 0x020E[31:0]  P0_DEN                      1                  0x00000001
-- 0x0212[47:0]  P1_NUM                      0                  0x000000000000
-- 0x0218[31:0]  P1_DEN                      0                  0x00000000
-- 0x021C[47:0]  P2_NUM                      0                  0x000000000000
-- 0x0222[31:0]  P2_DEN                      0                  0x00000000
-- 0x0226[47:0]  P3_NUM                      0                  0x000000000000
-- 0x022C[31:0]  P3_DEN                      0                  0x00000000
-- 0x0231[3:0]   P0_FRACN_MODE               11                 0xB
-- 0x0231[4]     P0_FRACN_EN                 0                  0x0
-- 0x0232[3:0]   P1_FRACN_MODE               11                 0xB
-- 0x0232[4]     P1_FRACN_EN                 0                  0x0
-- 0x0233[3:0]   P2_FRACN_MODE               11                 0xB
-- 0x0233[4]     P2_FRACN_EN                 0                  0x0
-- 0x0234[3:0]   P3_FRACN_MODE               11                 0xB
-- 0x0234[4]     P3_FRACN_EN                 0                  0x0
-- 0x0235[43:0]  MXAXB_NUM                   590558003200       0x08980000000
-- 0x023B[31:0]  MXAXB_DEN                   2147483648         0x80000000
-- 0x024A[23:0]  R0_REG                      0                  0x000000
-- 0x024D[23:0]  R1_REG                      0                  0x000000
-- 0x0250[23:0]  R2_REG                      0                  0x000000
-- 0x0253[23:0]  R3_REG                      0                  0x000000
-- 0x0256[23:0]  R4_REG                      0                  0x000000
-- 0x0259[23:0]  R5_REG                      0                  0x000000
-- 0x025C[23:0]  R6_REG                      0                  0x000000
-- 0x025F[23:0]  R7_REG                      0                  0x000000
-- 0x0262[23:0]  R8_REG                      0                  0x000000
-- 0x0268[23:0]  R9_REG                      0                  0x000000
-- 0x026B[7:0]   DESIGN_ID0                  115                0x73
-- 0x026C[7:0]   DESIGN_ID1                  80                 0x50
-- 0x026D[7:0]   DESIGN_ID2                  72                 0x48
-- 0x026E[7:0]   DESIGN_ID3                  88                 0x58
-- 0x026F[7:0]   DESIGN_ID4                  95                 0x5F
-- 0x0270[7:0]   DESIGN_ID5                  71                 0x47
-- 0x0271[7:0]   DESIGN_ID6                  84                 0x54
-- 0x0272[7:0]   DESIGN_ID7                  77                 0x4D
-- 0x028A[4:0]   OOF0_TRG_THR_EXT            0                  0x00
-- 0x028B[4:0]   OOF1_TRG_THR_EXT            0                  0x00
-- 0x028C[4:0]   OOF2_TRG_THR_EXT            0                  0x00
-- 0x028D[4:0]   OOF3_TRG_THR_EXT            0                  0x00
-- 0x028E[4:0]   OOF0_CLR_THR_EXT            0                  0x00
-- 0x028F[4:0]   OOF1_CLR_THR_EXT            0                  0x00
-- 0x0290[4:0]   OOF2_CLR_THR_EXT            0                  0x00
-- 0x0291[4:0]   OOF3_CLR_THR_EXT            0                  0x00
-- 0x0294[7:4]   FASTLOCK_EXTEND_SCL         11                 0xB
-- 0x0296[1]     LOL_SLW_VALWIN_SELX         1                  0x1
-- 0x0297[1]     FASTLOCK_DLY_ONSW_EN        1                  0x1
-- 0x0299[1]     FASTLOCK_DLY_ONLOL_EN       1                  0x1
-- 0x029D[19:0]  FASTLOCK_DLY_ONLOL          506                0x001FA
-- 0x02A9[19:0]  FASTLOCK_DLY_ONSW           1228               0x004CC
-- 0x02B7[3:2]   LOL_NOSIG_TIME              3                  0x3
-- 0x0302[43:0]  N0_NUM                      118111600640       0x01B80000000
-- 0x0308[31:0]  N0_DEN                      2147483648         0x80000000
-- 0x030C[0]     N0_UPDATE                   0                  0x0
-- 0x030D[43:0]  N1_NUM                      0                  0x00000000000
-- 0x0313[31:0]  N1_DEN                      0                  0x00000000
-- 0x0317[0]     N1_UPDATE                   0                  0x0
-- 0x0318[43:0]  N2_NUM                      0                  0x00000000000
-- 0x031E[31:0]  N2_DEN                      0                  0x00000000
-- 0x0322[0]     N2_UPDATE                   0                  0x0
-- 0x0323[43:0]  N3_NUM                      0                  0x00000000000
-- 0x0329[31:0]  N3_DEN                      0                  0x00000000
-- 0x032D[0]     N3_UPDATE                   0                  0x0
-- 0x032E[43:0]  N4_NUM                      0                  0x00000000000
-- 0x0334[31:0]  N4_DEN                      0                  0x00000000
-- 0x0338[0]     N4_UPDATE                   0                  0x0
-- 0x0338[1]     N_UPDATE                    0                  0x0
-- 0x0339[4:0]   N_FSTEP_MSK                 31                 0x1F
-- 0x033B[43:0]  N0_FSTEPW                   0                  0x00000000000
-- 0x0341[43:0]  N1_FSTEPW                   0                  0x00000000000
-- 0x0347[43:0]  N2_FSTEPW                   0                  0x00000000000
-- 0x034D[43:0]  N3_FSTEPW                   0                  0x00000000000
-- 0x0353[43:0]  N4_FSTEPW                   0                  0x00000000000
-- 0x0359[15:0]  N0_DELAY                    0                  0x0000
-- 0x035B[15:0]  N1_DELAY                    0                  0x0000
-- 0x035D[15:0]  N2_DELAY                    0                  0x0000
-- 0x035F[15:0]  N3_DELAY                    0                  0x0000
-- 0x0361[15:0]  N4_DELAY                    0                  0x0000
-- 0x0487[0]     ZDM_EN                      0                  0x0
-- 0x0487[2:1]   ZDM_IN_SEL                  0                  0x0
-- 0x0487[4]     ZDM_AUTOSW_EN               0                  0x0
-- 0x0508[5:0]   BW0_PLL                     19                 0x13
-- 0x0509[5:0]   BW1_PLL                     34                 0x22
-- 0x050A[5:0]   BW2_PLL                     12                 0x0C
-- 0x050B[5:0]   BW3_PLL                     11                 0x0B
-- 0x050C[5:0]   BW4_PLL                     7                  0x07
-- 0x050D[5:0]   BW5_PLL                     63                 0x3F
-- 0x050E[5:0]   FASTLOCK_BW0_PLL            22                 0x16
-- 0x050F[5:0]   FASTLOCK_BW1_PLL            42                 0x2A
-- 0x0510[5:0]   FASTLOCK_BW2_PLL            9                  0x09
-- 0x0511[5:0]   FASTLOCK_BW3_PLL            8                  0x08
-- 0x0512[5:0]   FASTLOCK_BW4_PLL            7                  0x07
-- 0x0513[5:0]   FASTLOCK_BW5_PLL            63                 0x3F
-- 0x0515[55:0]  M_NUM                       2834678415360      0x00029400000000
-- 0x051C[31:0]  M_DEN                       2147483648         0x80000000
-- 0x0521[3:0]   M_FRAC_MODE                 11                 0xB
-- 0x0521[4]     M_FRAC_EN                   0                  0x0
-- 0x0521[5]     PLL_OUT_RATE_SEL            1                  0x1
-- 0x052A[0]     IN_SEL_REGCTRL              1                  0x1
-- 0x052A[3:1]   IN_SEL                      0                  0x0
-- 0x052B[0]     FASTLOCK_AUTO_EN            1                  0x1
-- 0x052B[1]     FASTLOCK_MAN                0                  0x0
-- 0x052C[0]     HOLD_EN                     1                  0x1
-- 0x052C[3]     HOLD_RAMP_BYP               0                  0x0
-- 0x052C[4]     HOLDEXIT_BW_SEL1            0                  0x0
-- 0x052C[7:5]   RAMP_STEP_INTERVAL          4                  0x4
-- 0x052D[1]     HOLD_RAMPBYP_NOHIST         1                  0x1
-- 0x052E[4:0]   HOLD_HIST_LEN               25                 0x19
-- 0x052F[4:0]   HOLD_HIST_DELAY             25                 0x19
-- 0x0531[4:0]   HOLD_REF_COUNT_FRC          0                  0x00
-- 0x0532[23:0]  HOLD_15M_CYC_COUNT          834                0x000342
-- 0x0535[0]     FORCE_HOLD                  0                  0x0
-- 0x0536[1:0]   CLK_SWITCH_MODE             0                  0x0
-- 0x0536[2]     HSW_EN                      0                  0x0
-- 0x0537[3:0]   IN_LOS_MSK                  0                  0x0
-- 0x0537[7:4]   IN_OOF_MSK                  0                  0x0
-- 0x0538[2:0]   IN0_PRIORITY                0                  0x0
-- 0x0538[6:4]   IN1_PRIORITY                0                  0x0
-- 0x0539[2:0]   IN2_PRIORITY                0                  0x0
-- 0x0539[6:4]   IN3_PRIORITY                0                  0x0
-- 0x053A[1:0]   HSW_MODE                    2                  0x2
-- 0x053A[3:2]   HSW_PHMEAS_CTRL             0                  0x0
-- 0x053B[9:0]   HSW_PHMEAS_THR              3                  0x003
-- 0x053D[4:0]   HSW_COARSE_PM_LEN           17                 0x11
-- 0x053E[4:0]   HSW_COARSE_PM_DLY           6                  0x06
-- 0x0589[12:0]  CAP_SHORT_DELAY             13                 0x000D
-- 0x059B[1]     INIT_LP_CLOSE_HO            0                  0x0
-- 0x059B[4]     HOLD_PRESERVE_HIST          1                  0x1
-- 0x059B[5]     HOLD_FRZ_WITH_INTONLY       1                  0x1
-- 0x059B[6]     HOLDEXIT_BW_SEL0            1                  0x1
-- 0x059B[7]     HOLDEXIT_STD_BO             1                  0x1
-- 0x059D[5:0]   HOLDEXIT_BW0                19                 0x13
-- 0x059E[5:0]   HOLDEXIT_BW1                36                 0x24
-- 0x059F[5:0]   HOLDEXIT_BW2                12                 0x0C
-- 0x05A0[5:0]   HOLDEXIT_BW3                11                 0x0B
-- 0x05A1[5:0]   HOLDEXIT_BW4                7                  0x07
-- 0x05A2[5:0]   HOLDEXIT_BW5                63                 0x3F
-- 0x05A6[2:0]   RAMP_STEP_SIZE              3                  0x3
-- 0x05A6[3]     RAMP_SWITCH_EN              0                  0x0
-- 0x0802[15:0]  FIXREGSA0                   1333               0x0535
-- 0x0804[7:0]   FIXREGSD0                   0                  0x00
-- 0x0805[15:0]  FIXREGSA1                   0                  0x0000
-- 0x0807[7:0]   FIXREGSD1                   0                  0x00
-- 0x0808[15:0]  FIXREGSA2                   0                  0x0000
-- 0x080A[7:0]   FIXREGSD2                   0                  0x00
-- 0x080B[15:0]  FIXREGSA3                   0                  0x0000
-- 0x080D[7:0]   FIXREGSD3                   0                  0x00
-- 0x080E[15:0]  FIXREGSA4                   0                  0x0000
-- 0x0810[7:0]   FIXREGSD4                   0                  0x00
-- 0x0811[15:0]  FIXREGSA5                   0                  0x0000
-- 0x0813[7:0]   FIXREGSD5                   0                  0x00
-- 0x0814[15:0]  FIXREGSA6                   0                  0x0000
-- 0x0816[7:0]   FIXREGSD6                   0                  0x00
-- 0x0817[15:0]  FIXREGSA7                   0                  0x0000
-- 0x0819[7:0]   FIXREGSD7                   0                  0x00
-- 0x081A[15:0]  FIXREGSA8                   0                  0x0000
-- 0x081C[7:0]   FIXREGSD8                   0                  0x00
-- 0x081D[15:0]  FIXREGSA9                   0                  0x0000
-- 0x081F[7:0]   FIXREGSD9                   0                  0x00
-- 0x0820[15:0]  FIXREGSA10                  0                  0x0000
-- 0x0822[7:0]   FIXREGSD10                  0                  0x00
-- 0x0823[15:0]  FIXREGSA11                  0                  0x0000
-- 0x0825[7:0]   FIXREGSD11                  0                  0x00
-- 0x0826[15:0]  FIXREGSA12                  0                  0x0000
-- 0x0828[7:0]   FIXREGSD12                  0                  0x00
-- 0x0829[15:0]  FIXREGSA13                  0                  0x0000
-- 0x082B[7:0]   FIXREGSD13                  0                  0x00
-- 0x082C[15:0]  FIXREGSA14                  0                  0x0000
-- 0x082E[7:0]   FIXREGSD14                  0                  0x00
-- 0x082F[15:0]  FIXREGSA15                  0                  0x0000
-- 0x0831[7:0]   FIXREGSD15                  0                  0x00
-- 0x0832[15:0]  FIXREGSA16                  0                  0x0000
-- 0x0834[7:0]   FIXREGSD16                  0                  0x00
-- 0x0835[15:0]  FIXREGSA17                  0                  0x0000
-- 0x0837[7:0]   FIXREGSD17                  0                  0x00
-- 0x0838[15:0]  FIXREGSA18                  0                  0x0000
-- 0x083A[7:0]   FIXREGSD18                  0                  0x00
-- 0x083B[15:0]  FIXREGSA19                  0                  0x0000
-- 0x083D[7:0]   FIXREGSD19                  0                  0x00
-- 0x083E[15:0]  FIXREGSA20                  0                  0x0000
-- 0x0840[7:0]   FIXREGSD20                  0                  0x00
-- 0x0841[15:0]  FIXREGSA21                  0                  0x0000
-- 0x0843[7:0]   FIXREGSD21                  0                  0x00
-- 0x0844[15:0]  FIXREGSA22                  0                  0x0000
-- 0x0846[7:0]   FIXREGSD22                  0                  0x00
-- 0x0847[15:0]  FIXREGSA23                  0                  0x0000
-- 0x0849[7:0]   FIXREGSD23                  0                  0x00
-- 0x084A[15:0]  FIXREGSA24                  0                  0x0000
-- 0x084C[7:0]   FIXREGSD24                  0                  0x00
-- 0x084D[15:0]  FIXREGSA25                  0                  0x0000
-- 0x084F[7:0]   FIXREGSD25                  0                  0x00
-- 0x0850[15:0]  FIXREGSA26                  0                  0x0000
-- 0x0852[7:0]   FIXREGSD26                  0                  0x00
-- 0x0853[15:0]  FIXREGSA27                  0                  0x0000
-- 0x0855[7:0]   FIXREGSD27                  0                  0x00
-- 0x0856[15:0]  FIXREGSA28                  0                  0x0000
-- 0x0858[7:0]   FIXREGSD28                  0                  0x00
-- 0x0859[15:0]  FIXREGSA29                  0                  0x0000
-- 0x085B[7:0]   FIXREGSD29                  0                  0x00
-- 0x085C[15:0]  FIXREGSA30                  0                  0x0000
-- 0x085E[7:0]   FIXREGSD30                  0                  0x00
-- 0x085F[15:0]  FIXREGSA31                  0                  0x0000
-- 0x0861[7:0]   FIXREGSD31                  0                  0x00
-- 0x090E[0]     XAXB_EXTCLK_EN              0                  0x0
-- 0x0943[0]     IO_VDD_SEL                  0                  0x0
-- 0x0949[3:0]   IN_EN                       1                  0x1
-- 0x0949[7:4]   IN_PULSED_CMOS_EN           0                  0x0
-- 0x094A[3:0]   INX_TO_PFD_EN               1                  0x1
-- 0x094E[11:0]  REFCLK_HYS_SEL              585                0x249
-- 0x095E[0]     MXAXB_INTEGER               0                  0x0
-- 0x0A02[4:0]   N_ADD_0P5                   0                  0x00
-- 0x0A03[4:0]   N_CLK_TO_OUTX_EN            1                  0x01
-- 0x0A04[4:0]   N_PIBYP                     1                  0x01
-- 0x0A05[4:0]   N_PDNB                      1                  0x01
-- 0x0A14[3]     N0_HIGH_FREQ                0                  0x0
-- 0x0A1A[3]     N1_HIGH_FREQ                0                  0x0
-- 0x0A20[3]     N2_HIGH_FREQ                0                  0x0
-- 0x0A26[3]     N3_HIGH_FREQ                0                  0x0
-- 0x0A2C[3]     N4_HIGH_FREQ                0                  0x0
-- 0x0B44[3:0]   PDIV_FRACN_CLK_DIS          15                 0xF
-- 0x0B44[5]     FRACN_CLK_DIS_PLL           1                  0x1
-- 0x0B46[3:0]   LOS_CLK_DIS                 0                  0x0
-- 0x0B47[4:0]   OOF_CLK_DIS                 14                 0x0E
-- 0x0B48[4:0]   OOF_DIV_CLK_DIS             14                 0x0E
-- 0x0B4A[4:0]   N_CLK_DIS                   30                 0x1E
-- 0x0B57[11:0]  VCO_RESET_CALCODE           270                0x10E
-- 
-- 
-- 

end package si5345_register_pkg;
